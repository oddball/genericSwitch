`define   nbrOfPorts  2
`define   nbrOfBanks  4
`define   addresses   32
`define   serialWidth  8
`define   parrallelWidth 512
`define   nbrOfVirtualDestPort 32
